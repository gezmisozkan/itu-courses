/*
	150180005	Yağmur Çağlar
	
	150180010	Elif Arıkan
	
	150180059	Veysel Emre Köse
*/
//////////////////////////////////////////////-------------------------/////////////////////////////////////////////
//////////////////////////////////////////////GATE IMPLEMENTATION TESTS/////////////////////////////////////////////
//////////////////////////////////////////////-------------------------/////////////////////////////////////////////

module nand_test();
	reg i_1, i_2;
	
	wire o;
	
	nand_gate uut(.i_1(i_1), .i_2(i_2), .o(o));
	
	initial begin
		i_1=0; i_2=0; #250;
		i_1=1; i_2=0; #250;
		i_1=0; i_2=1; #250;
		i_1=1; i_2=1; #250;
	end
endmodule

//////////////////////////////////////////////-------------------------/////////////////////////////////////////////
//////////////////////////////////////////////-------PART 1 TESTS------/////////////////////////////////////////////
//////////////////////////////////////////////-------------------------/////////////////////////////////////////////

module sr_test();
	reg S, R;

	wire Q, Qnot;
	
	SR  uut(.S(S), .R(R), .Q(Q), .Qnot(Qnot));
	
	initial begin
		S=1; R=0; #200;
		S=0; R=0; #200;
		S=0; R=1; #200;
		S=0; R=0; #200;
		S=1; R=1; #200;
	end
endmodule

//////////////////////////////////////////////-------------------------/////////////////////////////////////////////
//////////////////////////////////////////////------PART 2 TEST--------/////////////////////////////////////////////
//////////////////////////////////////////////-------------------------/////////////////////////////////////////////
module sr_e_test();
	reg S, R,E;

	wire Q, Qnot;
	
	SR_E  uut(.S(S), .R(R), .E(E), .Q(Q), .Qnot(Qnot));
	
	initial begin
		S=0; E=0; R=0; #200;
		S=1; E=1; R=0; #200;
		S=0; E=1; R=1; #200;
		S=0; E=1; R=0; #200;
		S=1; E=1; R=1; #200; //forbidden
	end
endmodule

//////////////////////////////////////////////-------------------------/////////////////////////////////////////////
//////////////////////////////////////////////--------PART 3 TEST -----/////////////////////////////////////////////
//////////////////////////////////////////////-------------------------/////////////////////////////////////////////
module d_latch_test();
	reg D, Clk;

	wire Q, Qnot;
	
	d_latch  uut(.D(D), .Clk(Clk), .Q(Q), .Qnot(Qnot));
	
	initial begin
		D=0; Clk=0; #125;
		D=0; Clk=1; #125;
		D=1; Clk=0; #125;
		D=1; Clk=1; #125;
		D=0; Clk=0; #125;
		D=0; Clk=1; #125;
		D=1; Clk=0; #125;
		D=1; Clk=1; #125;
	end
endmodule


module d_flip_flop_test();
	reg D, Clk;

	wire Q, Qnot;
	
	d_flip_flop uut(.D(D), .Clk(Clk), .Q(Q), .Qnot(Qnot));
	
	initial begin
		D=0; Clk=0; #125;
		D=0; Clk=1; #125;
		D=1; Clk=0; #125;
		D=1; Clk=1; #125;
		D=0; Clk=0; #125;
		D=0; Clk=1; #125;
		D=1; Clk=0; #125;
		D=1; Clk=1; #125;
	end
endmodule

//////////////////////////////////////////////-------------------------/////////////////////////////////////////////
//////////////////////////////////////////////------PART 4 TEST -------/////////////////////////////////////////////
//////////////////////////////////////////////-------------------------/////////////////////////////////////////////

module part4_test();
       reg [15:0] yildik;
       reg clk;
       reg load;
       wire Q;
       
       shifreg uut(.yildik(yildik), .clk(clk), .load(load), .Q(Q));
       
       initial begin
            clk=0;
            yildik=16'b1010101010101010; load=1; #8;
            load=0; #128;
            yildik=16'b1100110011001100; load=1; #8;
            load=0; #128;
            yildik=16'b1111000011110000; load=1; #8;
            load=0; #128;
            yildik=16'b1000000010000000; load=1; #8;
            load=0; #128;
            yildik=16'b1000000000000000; load=1; #8;
            load=0; #128;
            yildik=16'b1110000000000000; load=1; #8;
            load=0; #128;
            yildik=16'b1111111111100000; load=1; #8;
            load=0; #128;
        end
        
        always begin 
            #4; clk=~clk;
        end 
endmodule 